//=======================================================
// register_renaming_unit.sv
//
// author: Woojin Jung
//=======================================================

import Type::*;

module RegRenamingUnit #(
  
)(
  input CLK,
  input RSTn,
  
  input Packet::DecoderToRru packetFromRru,
  
  output Packet::RruToRob1 packetToRob1,
  output Packet::RruToRob2 pacektToRob2
);
  
  
  
  
  
  
  
  
  
  
  
  
endmodule
